library ieee;
use ieee.std_logic_1164.all;
use ieee.Numeric_std.all;

entity riscy_vee is
	
	port(
			clk_50		: in std_logic
		);
	
	
end riscy_vee;

architecture desc of riscy_vee is

begin

end desc;
